module sawtooth_gen();


endmodule 